module sumaresta(

	input wire [1:0] A,
	input wire [3:0] Q,
	output wire [3:0] D
	);
	
	assign D[3] =
				(~A[1] & ~A[0] & Q[3]) | 
				(Q[3] & Q[1] & ~Q[0]) |
				(Q[3] & Q[2] & ~Q[1]) |
				(A[0] & Q[3] & ~Q[2]) |
				(A[1] & Q[3] & Q[0]) |
				(~A[1] & A[0] & ~Q[3] & Q[2] & Q[1] & Q[0]) |
				(A[1] & ~A[0] & ~Q[3] & ~Q[2] & ~Q[1] & ~Q[0]);
			
	assign D[2] =
				(~A[1] & ~A[0] & Q[2]) | 
				(Q[2] & Q[1] & ~Q[0]) |
				(A[0] & Q[2] & ~Q[1]) |
				(A[1] & Q[2] & Q[0]) |
				(~A[1] & A[0] & ~Q[2] & Q[1] & Q[0]) |
				(A[1] & ~A[0] & ~Q[2] & ~Q[1] & ~Q[0]);
			
	assign D[1] =
				(~A[1] & ~A[0] & Q[1])	| 
				(A[0] & Q[1] & ~Q[0])	|
				(A[1] & Q[1] & Q[0]) |
				(~A[1] & A[0] & ~Q[1] & Q[0]) |
				(A[1] & ~A[0] & ~Q[1] & ~Q[0]) ;
				
	assign D[0] =
				(~A[1] & ~A[0] & Q[0])	| 
				(~A[1] & A[0] & ~Q[0])	|
				(A[1] & ~A[0] & ~Q[0]) |
				(A[1] & A[0] & Q[0]) ;
			
	endmodule